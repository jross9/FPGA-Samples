// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		input  wire  clk_clk,       //   clk.clk
		output wire  hdmi_clk,      //  hdmi.clk
		input  wire  reset_reset_n,  // reset.reset_n
		output wire  reset_n
	);

	soc_system_pll_0 pll_0 (
		.refclk   (clk_clk),        //  refclk.clk
		.rst      (~reset_reset_n), //   reset.reset
		.outclk_0 (hdmi_clk),       // outclk0.clk
		.locked   (reset_n)         //  locked.export
	);

endmodule
